* Extracted by KLayout with SG13G2 LVS runset on : 23/06/2025 11:51

.SUBCKT inverter
M$1 \$1 \$4 \$3 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u
+ PD=1.34u
M$2 \$2 \$4 \$3 \$2 sg13_lv_pmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u
+ PD=1.34u
.ENDS inverter
