* Extracted by KLayout with SG13G2 LVS runset on : 18/06/2025 22:02

.SUBCKT TOP
M$1 \$2 \$5 \$3 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u
+ PD=1.34u
M$2 \$3 \$5 \$4 \$6 sg13_lv_pmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u
+ PD=1.34u
.ENDS TOP
