* Qucs 25.1.2  /home/mtfir/microelectronics/projects/ihp-inverter/qucs-s/inverter.sch
.INCLUDE "/usr/share/qucs-s/xspice_cmlib/include/ngspice_mathfunc.inc"

.SUBCKT IHP_PDK_nonlinear_components_sg13_lv_pmos gnd d g s b w=0.35u l=0.34u ng=1 m=1 mismatch=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346e-6 z2=0.38e-6 wmin=0.15e-6 rfmode=0 pre_layout=1 
X1 d g s b  sg13_lv_pmos w={w} l={l} ng={ng} m={1} mm_ok={mismatch} as={as} ad={ad} pd={pd} 
+ ps={ps} trise={trise} z1={z1} z2={z2} wmin={wmin} rfmode={rfmode} pre_layout={pre_layout}
.ENDS
  

.SUBCKT IHP_PDK_nonlinear_components_sg13_lv_nmos gnd d g s b w=0.35u l=0.34u ng=1 m=1 mismatch=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346e-6 z2=0.38e-6 wmin=0.15e-6 rfmode=0 pre_layout=1 mlist=1
X1 d g s b  sg13_lv_nmos w={w} l={l} ng={ng} m={m} mm_ok={mismatch} as={as} ad={ad} pd={pd} 
+ ps={ps} trise={trise} z1={z1} z2={z2} wmin={wmin} rfmode={rfmode} pre_layout={pre_layout}
.ENDS
  
.LIB cornerMOSlv.lib mos_tt

Xsg13_lv_pmos1 0  VCC VIN _net0 VOUT IHP_PDK_nonlinear_components_sg13_lv_pmos w=0.35U l=0.34U ng=1 m=1 mismatch=0 as=0 ad=0 pd=0 ps=0 trise=0.346E-6 z1=0.38E-6 z2=0.15E-6 wmin=0 rfmode=1 pre_layout=1
Xsg13_lv_nmos1 0  _net0 VIN VDD VOUT IHP_PDK_nonlinear_components_sg13_lv_nmos w=0.35U l=0.34U ng=1 m=1 mismatch=0 as=0 ad=0 pd=0 ps=0 trise=0.346E-6 z1=0.38E-6 z2=0.15E-6 wmin=0 rfmode=1 pre_layout=1


.control

exit
.endc
.END
