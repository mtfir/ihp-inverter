** sch_path: /home/mtfir/microelectronics/projects/ihp-inverter/xschem/inverter.sch
.SUBCKT inverter A Y VDD VSS
*.PININFO A:I Y:O VDD:B VSS:B
M1 Y A VSS VSS sg13_lv_nmos w=150n l=130n ng=1 m=1
M2 Y A VDD VDD sg13_lv_pmos w=150n l=130n ng=1 m=1
.ENDS
