** sch_path: /home/mtfir/microelectronics/projects/ihp-inverter/xschem/inverter.sch
**.subckt inverter A Y VDD VSS
*.ipin A
*.opin Y
*.iopin VDD
*.iopin VSS
XM1 Y A VSS VSS sg13_lv_nmos w=150n l=130n ng=1 m=1 rfmode=1
XM2 Y A VDD VDD sg13_lv_pmos w=150n l=130n ng=1 m=1 rfmode=1
**.ends
.end
